/*
 * constants.vh
 *
 * Definitions for commonly used constants.
 */

`ifndef _constants_vh
`define _constants_vh

localparam  BIT_WIDTH = 32;

`endif