/*
 * constants.vh
 *
 * Definitions for commonly used constants.
 */

`ifndef _constants_vh
`define _constants_vh

package constants;
    localparam  REGFILE_SIZE = 32;
    localparam  WORD_LENGTH = 32;
endpackage;

`endif